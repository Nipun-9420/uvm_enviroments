    /*
    only basic output with configuration for nu of agent 
    --------------------------------------------------------------
Name                       Type                    Size  Value
--------------------------------------------------------------
uvm_test_top               router_test             -     @336 
  dst_agtt                 dst_agent_top           -     @349 
    dst_agh[0]             dst_agent               -     @374 
      ddrvh                dst_driver              -     @465 
        rsp_port           uvm_analysis_port       -     @484 
        seq_item_port      uvm_seq_item_pull_port  -     @474 
      dmonh                dst_monitor             -     @494 
      dseqrh               dst_sequencer           -     @503 
        rsp_export         uvm_analysis_export     -     @512 
        seq_item_export    uvm_seq_item_pull_imp   -     @630 
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    dst_agh[1]             dst_agent               -     @383 
      ddrvh                dst_driver              -     @646 
        rsp_port           uvm_analysis_port       -     @665 
        seq_item_port      uvm_seq_item_pull_port  -     @655 
      dmonh                dst_monitor             -     @675 
      dseqrh               dst_sequencer           -     @684 
        rsp_export         uvm_analysis_export     -     @693 
        seq_item_export    uvm_seq_item_pull_imp   -     @811 
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    dst_agh[2]             dst_agent               -     @392 
      ddrvh                dst_driver              -     @827 
        rsp_port           uvm_analysis_port       -     @846 
        seq_item_port      uvm_seq_item_pull_port  -     @836 
      dmonh                dst_monitor             -     @856 
      dseqrh               dst_sequencer           -     @865 
        rsp_export         uvm_analysis_export     -     @874 
        seq_item_export    uvm_seq_item_pull_imp   -     @992 
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    dst_agh[3]             dst_agent               -     @401 
      ddrvh                dst_driver              -     @1008
        rsp_port           uvm_analysis_port       -     @1027
        seq_item_port      uvm_seq_item_pull_port  -     @1017
      dmonh                dst_monitor             -     @1037
      dseqrh               dst_sequencer           -     @1046
        rsp_export         uvm_analysis_export     -     @1055
        seq_item_export    uvm_seq_item_pull_imp   -     @1173
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    dst_agh[4]             dst_agent               -     @410 
      ddrvh                dst_driver              -     @1189
        rsp_port           uvm_analysis_port       -     @1208
        seq_item_port      uvm_seq_item_pull_port  -     @1198
      dmonh                dst_monitor             -     @1218
      dseqrh               dst_sequencer           -     @1227
        rsp_export         uvm_analysis_export     -     @1236
        seq_item_export    uvm_seq_item_pull_imp   -     @1354
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    dst_agh[5]             dst_agent               -     @419 
      ddrvh                dst_driver              -     @1370
        rsp_port           uvm_analysis_port       -     @1389
        seq_item_port      uvm_seq_item_pull_port  -     @1379
      dmonh                dst_monitor             -     @1399
      dseqrh               dst_sequencer           -     @1408
        rsp_export         uvm_analysis_export     -     @1417
        seq_item_export    uvm_seq_item_pull_imp   -     @1535
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    dst_agh[6]             dst_agent               -     @428 
      ddrvh                dst_driver              -     @1551
        rsp_port           uvm_analysis_port       -     @1570
        seq_item_port      uvm_seq_item_pull_port  -     @1560
      dmonh                dst_monitor             -     @1580
      dseqrh               dst_sequencer           -     @1589
        rsp_export         uvm_analysis_export     -     @1598
        seq_item_export    uvm_seq_item_pull_imp   -     @1716
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    dst_agh[7]             dst_agent               -     @437 
      ddrvh                dst_driver              -     @1732
        rsp_port           uvm_analysis_port       -     @1751
        seq_item_port      uvm_seq_item_pull_port  -     @1741
      dmonh                dst_monitor             -     @1761
      dseqrh               dst_sequencer           -     @1770
        rsp_export         uvm_analysis_export     -     @1779
        seq_item_export    uvm_seq_item_pull_imp   -     @1897
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    dst_agh[8]             dst_agent               -     @446 
      ddrvh                dst_driver              -     @1913
        rsp_port           uvm_analysis_port       -     @1932
        seq_item_port      uvm_seq_item_pull_port  -     @1922
      dmonh                dst_monitor             -     @1942
      dseqrh               dst_sequencer           -     @1951
        rsp_export         uvm_analysis_export     -     @1960
        seq_item_export    uvm_seq_item_pull_imp   -     @2078
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    dst_agh[9]             dst_agent               -     @455 
      ddrvh                dst_driver              -     @2094
        rsp_port           uvm_analysis_port       -     @2113
        seq_item_port      uvm_seq_item_pull_port  -     @2103
      dmonh                dst_monitor             -     @2123
      dseqrh               dst_sequencer           -     @2132
        rsp_export         uvm_analysis_export     -     @2141
        seq_item_export    uvm_seq_item_pull_imp   -     @2259
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
  src_agtt                 src_agent_top           -     @358 
    src_agh[0]             src_agent               -     @2275
      sdrvh                src_driver              -     @2339
        rsp_port           uvm_analysis_port       -     @2358
        seq_item_port      uvm_seq_item_pull_port  -     @2348
      smonh                src_monitor             -     @2368
      sseqrh               src_sequencer           -     @2377
        rsp_export         uvm_analysis_export     -     @2386
        seq_item_export    uvm_seq_item_pull_imp   -     @2504
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    src_agh[1]             src_agent               -     @2284
      sdrvh                src_driver              -     @2520
        rsp_port           uvm_analysis_port       -     @2539
        seq_item_port      uvm_seq_item_pull_port  -     @2529
      smonh                src_monitor             -     @2549
      sseqrh               src_sequencer           -     @2558
        rsp_export         uvm_analysis_export     -     @2567
        seq_item_export    uvm_seq_item_pull_imp   -     @2685
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    src_agh[2]             src_agent               -     @2293
      sdrvh                src_driver              -     @2701
        rsp_port           uvm_analysis_port       -     @2720
        seq_item_port      uvm_seq_item_pull_port  -     @2710
      smonh                src_monitor             -     @2730
      sseqrh               src_sequencer           -     @2739
        rsp_export         uvm_analysis_export     -     @2748
        seq_item_export    uvm_seq_item_pull_imp   -     @2866
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    src_agh[3]             src_agent               -     @2302
      sdrvh                src_driver              -     @2882
        rsp_port           uvm_analysis_port       -     @2901
        seq_item_port      uvm_seq_item_pull_port  -     @2891
      smonh                src_monitor             -     @2911
      sseqrh               src_sequencer           -     @2920
        rsp_export         uvm_analysis_export     -     @2929
        seq_item_export    uvm_seq_item_pull_imp   -     @3047
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    src_agh[4]             src_agent               -     @2311
      sdrvh                src_driver              -     @3063
        rsp_port           uvm_analysis_port       -     @3082
        seq_item_port      uvm_seq_item_pull_port  -     @3072
      smonh                src_monitor             -     @3092
      sseqrh               src_sequencer           -     @3101
        rsp_export         uvm_analysis_export     -     @3110
        seq_item_export    uvm_seq_item_pull_imp   -     @3228
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    src_agh[5]             src_agent               -     @2320
      sdrvh                src_driver              -     @3244
        rsp_port           uvm_analysis_port       -     @3263
        seq_item_port      uvm_seq_item_pull_port  -     @3253
      smonh                src_monitor             -     @3273
      sseqrh               src_sequencer           -     @3282
        rsp_export         uvm_analysis_export     -     @3291
        seq_item_export    uvm_seq_item_pull_imp   -     @3409
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
    src_agh[6]             src_agent               -     @2329
      sdrvh                src_driver              -     @3425
        rsp_port           uvm_analysis_port       -     @3444
        seq_item_port      uvm_seq_item_pull_port  -     @3434
      smonh                src_monitor             -     @3454
      sseqrh               src_sequencer           -     @3463
        rsp_export         uvm_analysis_export     -     @3472
        seq_item_export    uvm_seq_item_pull_imp   -     @3590
        arbitration_queue  array                   0     -    
        lock_queue         array                   0     -    
        num_last_reqs      integral                32    'd1  
        num_last_rsps      integral                32    'd1  
--------------------------------------------------------------

    */

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    typedef enum {UVM_ACTIVE,UVM_PASSIVE} uvm_active_passive_enum;

    //#################################################################################  SORCE

    //================================
    //================================   XTN
    //================================

    class src_config extends uvm_object;
        `uvm_object_utils(src_config)

        function new(string name ="src_config");
                super.new(name);
        endfunction

    endclass
    class src_xtn extends uvm_sequence_item;
        `uvm_object_utils(src_xtn)
        function new(string name ="src_xtn");
            super.new(name);
        endfunction //new()
    endclass 


    //================================
    //================================   sequence
    //================================
    class src_seq extends uvm_sequence #(src_xtn);
        `uvm_object_utils(src_seq)
        function new(string name ="src_seq");
            super.new(name);
        endfunction //new()
    endclass //src_seq extends superClass


    //================================
    //================================   monitor
    //================================
    class src_monitor extends uvm_monitor;
        `uvm_component_utils(src_monitor)
        function new(string name ="src_monitor",uvm_component parent);
            super.new(name,parent);
        endfunction //new()
    endclass //src_monitor extends superClass


    //================================
    //================================   driver
    //================================
    class src_driver extends uvm_driver #(src_xtn);
        `uvm_component_utils(src_driver)
        function new(string name ="src_driver",uvm_component parent);
            super.new(name,parent);
        endfunction //new()
    endclass //src_driver



    //================================
    //================================   sequencer
    //================================
    class src_sequencer extends uvm_sequencer #(src_xtn);
        `uvm_component_utils(src_sequencer)
        function new(string name ="src_sequencer",uvm_component parent);
            super.new(name,parent);
        endfunction //new()
    endclass //src_driver

    //================================
    //================================   src_agent
    //================================
    class src_agent extends uvm_agent;
        `uvm_component_utils(src_agent)
        src_driver     sdrvh;
        src_monitor    smonh;
        src_sequencer sseqrh;
        function new(string name ="src_agent",uvm_component parent);
            super.new(name,parent);
        endfunction //new()

        function void build_phase(uvm_phase phase);
            super.build_phase(phase);
            sdrvh = src_driver::type_id::create("sdrvh",this);
            smonh = src_monitor::type_id::create("smonh",this);
            sseqrh = src_sequencer::type_id::create("sseqrh",this);
        endfunction
    endclass //src_agent extends superClass


    //================================
    //================================   src_agent_top
    //================================
    class src_agent_top extends uvm_env;
        `uvm_component_utils(src_agent_top)
        int no_src_agent;
        src_agent src_agh[];
        function new(string name ="src_agent_top",uvm_component parent);
            super.new(name,parent);
        endfunction //new()

        function void build_phase(uvm_phase phase);
            super.build_phase(phase);

            if(! uvm_config_db#(int)::get(this, "", "no_src_agent", no_src_agent))
            `uvm_fatal(get_name(), "failinf no of dst agt")
            
            src_agh = new[no_src_agent];
            foreach (src_agh[i]) 
            begin
                src_agh[i] = src_agent::type_id::create($sformatf("src_agh[%0d]",i),this);
            end

        endfunction
    endclass //src_agent extends superClass






    //#################################################################################  DESTINATION


    class dst_xtn extends uvm_sequence_item;
        `uvm_object_utils(dst_xtn)
        function new(string name ="dst_xtn");
            super.new(name);
        endfunction //new()
    endclass 


    //================================
    //================================   sequence
    //================================
    class dst_seq extends uvm_sequence #(dst_xtn);
        `uvm_object_utils(dst_seq)
        function new(string name ="dst_seq");
            super.new(name);
        endfunction //new()
    endclass //dst_seq extends superClass


    //================================
    //================================   monitor
    //================================
    class dst_monitor extends uvm_monitor;
        `uvm_component_utils(dst_monitor)
        
        function new(string name ="dst_monitor",uvm_component parent);
            super.new(name,parent);
        endfunction //new()
    endclass //dst_monitor extends superClass


    //================================
    //================================   driver
    //================================
    class dst_driver extends uvm_driver #(dst_xtn);
        `uvm_component_utils(dst_driver)
        function new(string name ="dst_driver",uvm_component parent);
            super.new(name,parent);
        endfunction //new()
    endclass //dst_driver



    //================================
    //================================   sequencer
    //================================
    class dst_sequencer extends uvm_sequencer#(dst_xtn);
        `uvm_component_utils(dst_sequencer)
        function new(string name ="dst_sequencer",uvm_component parent);
            super.new(name,parent);
        endfunction //new()
    endclass //dst_driver


    //================================
    //================================   dst_agent
    //================================
    class dst_agent extends uvm_agent;
        `uvm_component_utils(dst_agent)

        dst_driver     ddrvh;
        dst_monitor    dmonh;
        dst_sequencer dseqrh;
        function new(string name ="dst_agent",uvm_component parent);
            super.new(name,parent);
        endfunction //new()

        function void build_phase(uvm_phase phase);
            super.build_phase(phase);
            ddrvh = dst_driver::type_id::create("ddrvh",this);
            dmonh = dst_monitor::type_id::create("dmonh",this);
            dseqrh = dst_sequencer::type_id::create("dseqrh",this);
        endfunction
    endclass //dst_agent extends superClass


    //================================
    //================================   ----------------------------------------------------------dst_agent_top
    //================================
    class dst_agent_top extends uvm_env;
        `uvm_component_utils(dst_agent_top)
        int no_dst_agent ;

        dst_agent dst_agh[];
        function new(string name ="dst_agent_top",uvm_component parent);
            super.new(name,parent);
        endfunction //new()

        function void build_phase(uvm_phase phase);
            super.build_phase(phase);
        if(! uvm_config_db#(int)::get(this, "", "no_dst_agent", no_dst_agent))
            `uvm_fatal(get_name(), "failinf no of dst agt")
            
            dst_agh = new[no_dst_agent];
            foreach (dst_agh[i]) 
            begin
                dst_agh[i] = dst_agent::type_id::create($sformatf("dst_agh[%0d]",i),this);
            end
                    
        endfunction

        function void end_of_elaboration_phase(uvm_phase phase);
            super.end_of_elaboration_phase(phase);
            uvm_top.print_topology();
        endfunction

    endclass //dst_agent extends superClass









    //#################################################################################  enviroment


    class route_env extends uvm_env;
        `uvm_component_utils(route_env)

        dst_agent_top dst_agtt;
        src_agent_top src_agtt;
        function new(string name ="route_env",uvm_component parent);
            super.new(name,parent);
        endfunction //new()

        function void build_phase(uvm_phase phase);
            super.build_phase(phase);
            dst_agtt = dst_agent_top::type_id::create("dst_agtt",this);
            src_agtt = src_agent_top::type_id::create("src_agtt",this);
        endfunction

        
        
    endclass //dst_agent extends superClass

    //#################################################################################  enviroment


    class router_test extends uvm_test;
        `uvm_component_utils(router_test)
        int no_src_agent =7;
        int no_dst_agent =10;
        dst_agent_top dst_agtt;
        src_agent_top src_agtt;
        function new(string name ="route_env",uvm_component parent);
            super.new(name,parent);
        endfunction //new()

        function void build_phase(uvm_phase phase);
            super.build_phase(phase);
            dst_agtt = dst_agent_top::type_id::create("dst_agtt",this);
            src_agtt = src_agent_top::type_id::create("src_agtt",this);

            uvm_config_db#(int)::set(this, "*", "no_src_agent", no_src_agent);
            uvm_config_db#(int)::set(this, "*", "no_dst_agent", no_dst_agent);
        endfunction
    endclass //dst_agent extends superClass


    module top; 
        initial 
            run_test("router_test");
        
        
    endmodule